`ifndef APB_PKG_SV
`define APB_PKG_SV
package ApbPkg;
//-------------------------------------------------------
//define
//-------------------------------------------------------
// `define TEST_TOP top

//-------------------------------------------------------
//parameter
//-------------------------------------------------------
localparam APB_DW  = 32;
localparam APB_AW  = 32;

//-------------------------------------------------------
//function
//-------------------------------------------------------

//-------------------------------------------------------
//task
//-------------------------------------------------------

endpackage
`endif //APB_PKG_SV
