//1.function define--------------------------
//2.report define-----------------------------
//3.implement define--------------------------


//#1.function define
`define COM_SYNC_STAGE      3
`define COM_MCFG_W          4

//#2.report define
`define COM_REPORT_ON
`define COM_ASSERT_ON

//#3.implement define
`define COM_RAM_AS_REG
`define COM_CDC_AS_REG
`define COM_CLKGATE_AS_LATCH

//`define COM_FPGA